`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Team Members:
// Overall percent effort of each team member:
// Brett Bushnell -- 50%
// Derek Mcmullen -- 50% 
// 
////////////////////////////////////////////////////////////////////////////////

module WriteBackUnit(RegWriteIn, MemToRegIn, ALUIn, MemoryReadDataIn, DestinationRegIn, RegWriteOut, RegWriteDataOut, DestinationRegOut);
	
    /* Control Signals*/
    output RegWriteOut; 
    /* Data Signals*/
    output [31:0] RegWriteDataOut;
    output [4:0] DestinationRegOut; 
	
	/* Control Signals*/
    input RegWriteIn; 
    input MemToRegIn; 
    /* Data Signals*/
    input [31:0] ALUIn;
    input [31:0] MemoryReadDataIn; 
    input [4:0] DestinationRegIn; 
    
    // Included Modules
	Mux32Bit2To1 Mux32Bit2To1_1(RegWriteDataOut, MemoryReadDataIn, ALUIn, MemToRegIn); 
	// TODO: need output mux for write data to mux in the JAL info to $RA(31)
	// TODO: need output mux for writeregister to hardwire in an option for $RA(31) 5 bits
	// should be controlled by 2 bits of jump or'd together
	
	// Assign statements
	assign RegWriteOut = RegWriteIn; 
	assign DestinationRegOut = DestinationRegIn;
    
endmodule

