`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Team Members:
// Overall percent effort of each team member:
// Brett Bushnell -- 50%
// Derek Mcmullen -- 50% 
//
////////////////////////////////////////////////////////////////////////////////

module Controller(Instruction, Branch, MemRead, MemWrite, RegWrite, MemToReg, RegDst, ALUOp, ALUSrc, HiLoALUControl, AddToHi, AddToLo, MoveToHi, HiLoSel, ZeroExtend, AltALUSrc1, ZeroALUSrc1, ZeroALUSrc2, Swap, ALUHiLoSelect, MOVN, MOVZ, StraightToHi, StraightToLo, LoadStoreByte, LoadStoreHalf, NotZero, Jump);
    
    /* Control Signals*/
    output reg Branch; 
    output reg MemRead; 
    output reg MemWrite; 
    output reg RegWrite; 
    output reg MemToReg; 
    output reg RegDst; 
    output reg [4:0] ALUOp; 
    output reg ALUSrc;
    output reg HiLoALUControl, AddToHi, AddToLo, MoveToHi, HiLoSel;
    output reg ZeroExtend; 
    output reg AltALUSrc1;
    output reg ZeroALUSrc1;
    output reg ZeroALUSrc2;
    output reg Swap; 
    output reg ALUHiLoSelect; 
    output reg MOVN;
    output reg MOVZ;
    output reg StraightToHi; 
    output reg StraightToLo;
    output reg LoadStoreByte;
    output reg LoadStoreHalf;
    output reg NotZero;
    output reg [1:0] Jump; 

    
    input [31:0] Instruction; 
    
    initial begin
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'bxxxxx;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0; 
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
    end


    // Decode the Instruction
    always @(Instruction) begin
    
    casex (Instruction)
     32'b00000000000000000000000000000000:    begin   // NOP Command
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'bXXXXX;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    
    /* ARITHMETIC OPS */
     32'b000000xxxxxxxxxxxxxxxxxxxx100000:    begin    // ADD Command
        RegWrite        <= 1'b1; 
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00010;
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
     32'b001001xxxxxxxxxxxxxxxxxxxxxxxxxx:    begin   // ADDIU Command
        RegWrite        <= 1'b1; 
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b00010;
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
     32'b000000xxxxxxxxxxxxxxxxxxxx100001:    begin   // ADDU Command
        RegWrite        <= 1'b1; 
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00010;
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
     32'b001000xxxxxxxxxxxxxxxxxxxxxxxxxx:    begin   // ADDI Command
        RegWrite        <= 1'b1; 
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b00010;
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
     32'b000000xxxxxxxxxxxxxxxxxxxx100010:    begin   // SUB Command
        RegWrite        <= 1'b1; 
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00110;
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0;
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
     32'b011100xxxxxxxxxxxxxxxxxxxx000010:    begin   // MUL Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b01000;
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
     32'b000000xxxxxxxxxxxxxxxxxxxx011000:    begin   // MULT Command
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b01000;
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b1; 
        StraightToLo    <= 1'b1;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
     32'b000000xxxxxxxxxxxxxxxxxxxx011001:    begin   // MULTU Command
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b10001;
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b1; 
        StraightToLo    <= 1'b1;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
     32'b011100xxxxxxxxxxxxxxxxxxxx000000:    begin   // MADD Command
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b01000;
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b1; 
        AddToLo         <= 1'b1; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
     32'b011100xxxxxxxxxxxxxxxxxxxx000100:    begin   // MSUB Command
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b01000;
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b1; 
        AddToHi         <= 1'b1; 
        AddToLo         <= 1'b1; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end   
      
    /* LOGICAL OPS*/
    32'b000000xxxxxxxxxxxxxxxxxxxx100100:    begin   // AND Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00000;
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b001100xxxxxxxxxxxxxxxxxxxxxxxxxx:    begin   // ANDI Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b00000;
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b1; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end   
    32'b000000xxxxxxxxxxxxxxxxxxxx100101:    begin   // OR Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00001;
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
     32'b000000xxxxxxxxxxxxxxxxxxxx100111:    begin   // NOR Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00011;
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0;  
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end   
    32'b000000xxxxxxxxxxxxxxxxxxxx100110:    begin   // XOR Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00100;
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b001101xxxxxxxxxxxxxxxxxxxxxxxxxx:    begin   // ORI Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b00001;
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b1; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0;
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end        
    32'b001110xxxxxxxxxxxxxxxxxxxxxxxxxx:    begin   // XORI Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b00100;       //need XOR
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b01111100000xxxxxxxxxx11000100000:    begin   // SEH Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b01001;       //need SEH
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end   
    32'b000000xxxxxxxxxxxxxxxxxxxx000000:    begin   // SLL Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b01011;      //need SLL
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b1; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b00000000000xxxxxxxxxxxxxxx000010:    begin   // SRL Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b01100;      //need SRL
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b1; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end  
    32'b000000xxxxxxxxxxxxxxxxxxxx000100:    begin   // SLLV Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00101;     //need SLLV
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b1; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b000000xxxxxxxxxxxxxxx00000000110:    begin   // SRLV Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b01111;     //need SRL
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b1; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end     
    32'b000000xxxxxxxxxxxxxxxxxxxx101010:    begin   // SLT Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00111;    
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b001010xxxxxxxxxxxxxxxxxxxxxxxxxx:    begin   // SLTI Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b00111;     
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b000000xxxxxxxxxxxxxxxxxxxx001011:    begin   // MOVN Command
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00010;     // need ADD
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b1;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b1;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b000000xxxxxxxxxxxxxxxxxxxx001010:    begin   // MOVZ Command
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00010;     // need ADD
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b1;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b1;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end     
    32'b000000xxxxxxxxxxxxxxx00001000110:    begin   // ROTRV Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b10000;     //need ROTRV
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b1; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0; 
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b00000000001xxxxxxxxxxxxxxx000010:    begin   // ROTR Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b01101;     //need ROTR
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b1; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b000000xxxxxxxxxxxxxxxxxxxx000011:    begin   // SRA Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b01110;     //need SRA
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b1; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b000000xxxxxxxxxxxxxxxxxxxx000111:    begin   // SRAV Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b01110;     //need SRA
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b1; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end    
    32'b01111100000xxxxxxxxxx10000100000:    begin   // SEB Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b01010;     //need SEB
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b001011xxxxxxxxxxxxxxxxxxxxxxxxxx:    begin   // SLTIU Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b10010;     //SLTU   
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end      
    32'b000000xxxxxxxxxxxxxxxxxxxx101011:    begin   // SLTU Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b10010;        //SLTU 
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;  
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b000000xxxxxxxxxxxxxxxxxxxx010001:    begin   // MTHI Command
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00010;        //ADD 
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b1;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b1; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0; 
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b000000xxxxxxxxxxxxxxxxxxxx010011:    begin   // MTLO Command
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00010;        //ADD 
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b1;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b1; 
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end 
    32'b0000000000000000xxxxx00000010000:    begin   // MFHI Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00010;        //ADD 
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b1;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b1; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0; 
        HiLoSel         <= 1'b1; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end                 
    32'b0000000000000000xxxxx00000010010:    begin   // MFLO Command
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00010;        //ADD 
        RegDst          <= 1'b1; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b1;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b1; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0; 
        HiLoSel         <= 1'b0; 
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b100011xxxxxxxxxxxxxxxxxxxxxxxxxx:   begin //LW
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b00010;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b1; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
    end
    32'b101011xxxxxxxxxxxxxxxxxxxxxxxxxx:   begin //SW
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b00010;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b1; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
    end
    32'b101000xxxxxxxxxxxxxxxxxxxxxxxxxx:   begin //SB
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b00010;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b1; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b1;
        LoadStoreHalf   <= 1'b0;
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
    end      
    32'b100001xxxxxxxxxxxxxxxxxxxxxxxxxx:   begin //LH
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b00010;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b1; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b1;
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
    end
    32'b100000xxxxxxxxxxxxxxxxxxxxxxxxxx:   begin //LB
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b00010;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b1; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b1;
        LoadStoreHalf   <= 1'b0;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b101001xxxxxxxxxxxxxxxxxxxxxxxxxx:   begin //SH
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b00010;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b1; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0; 
        ZeroALUSrc2     <= 1'b0;
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b1;      
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end
    32'b00111100000xxxxxxxxxxxxxxxxxxxxx:   begin //LUI
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b1;
        ALUOp           <= 5'b10011;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b1; 
        MemToReg        <= 1'b1;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0;    
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
      end

    32'b000001xxxxx00001xxxxxxxxxxxxxxxx:   begin //BGEZ
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b10100;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b1; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b1; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0; 
        NotZero         <= 1'b1;
        Jump            <= 2'b00;
    end

    32'b000100xxxxxxxxxxxxxxxxxxxxxxxxxx:   begin // BEQ
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00100;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b1; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0; 
        NotZero         <= 1'b0;
        Jump            <= 2'b00;
    end

    32'b000101xxxxxxxxxxxxxxxxxxxxxxxxxx:   begin // BNE
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00100;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b1; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0; 
        NotZero         <= 1'b1;
        Jump            <= 2'b00;
    end

    32'b000111xxxxx00000xxxxxxxxxxxxxxxx:   begin // BGTZ
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00111;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b1; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b1; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0; 
        NotZero         <= 1'b1;
        Jump            <= 2'b00;
    end

    32'b000110xxxxx00000xxxxxxxxxxxxxxxx:   begin // BLEZ
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b10100;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b1; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b1; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0; 
        NotZero         <= 1'b1;
        Jump            <= 2'b00;
    end

    32'b000001xxxxx00000xxxxxxxxxxxxxxxx:   begin // BLTZ
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'b00111;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b1; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0; 
        NotZero         <= 1'b1;
        Jump            <= 2'b00;
    end
    
    32'b000010xxxxxxxxxxxxxxxxxxxxxxxxxx:   begin // J
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'bXXXXX;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0; 
        NotZero         <= 1'b0;
        Jump            <= 2'b01;
    end    

    32'b000000xxxxx0000000000xxxxx001000:   begin // JR
        RegWrite        <= 1'b0;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'bXXXXX;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0; 
        NotZero         <= 1'b0;
        Jump            <= 2'b10;
    end     

    32'b000011xxxxxxxxxxxxxxxxxxxxxxxxxx:   begin // JAL
        RegWrite        <= 1'b1;
        ALUSrc          <= 1'b0;
        ALUOp           <= 5'bXXXXX;        
        RegDst          <= 1'b0; 
        Branch          <= 1'b0; 
        MemWrite        <= 1'b0; 
        MemRead         <= 1'b0; 
        ZeroExtend      <= 1'b0; 
        MemToReg        <= 1'b0;
        AltALUSrc1      <= 1'b0; 
        ZeroALUSrc1     <= 1'b0;
        ZeroALUSrc2     <= 1'b0; 
        Swap            <= 1'b0; 
        ALUHiLoSelect   <= 1'b0; 
        HiLoALUControl  <= 1'b0; 
        AddToHi         <= 1'b0; 
        AddToLo         <= 1'b0; 
        MoveToHi        <= 1'b0; 
        StraightToHi    <= 1'b0; 
        StraightToLo    <= 1'b0;
        HiLoSel         <= 1'b0;
        MOVN            <= 1'b0;
        MOVZ            <= 1'b0;
        LoadStoreByte   <= 1'b0;
        LoadStoreHalf   <= 1'b0; 
        NotZero         <= 1'b0;
        Jump            <= 2'b01;
    end
    default: begin
        RegWrite        <= 1'b0;
            ALUSrc          <= 1'b0;
            ALUOp           <= 5'b00000;        
            RegDst          <= 1'b0; 
            Branch          <= 1'b0; 
            MemWrite        <= 1'b0; 
            MemRead         <= 1'b0; 
            ZeroExtend      <= 1'b0; 
            MemToReg        <= 1'b0;
            AltALUSrc1      <= 1'b0; 
            ZeroALUSrc1     <= 1'b0;
            ZeroALUSrc2     <= 1'b0; 
            Swap            <= 1'b0; 
            ALUHiLoSelect   <= 1'b0; 
            HiLoALUControl  <= 1'b0; 
            AddToHi         <= 1'b0; 
            AddToLo         <= 1'b0; 
            MoveToHi        <= 1'b0; 
            StraightToHi    <= 1'b0; 
            StraightToLo    <= 1'b0;
            HiLoSel         <= 1'b0;
            MOVN            <= 1'b0;
            MOVZ            <= 1'b0;
            LoadStoreByte   <= 1'b0;
            LoadStoreHalf   <= 1'b0; 
            NotZero         <= 1'b0;
            Jump            <= 2'b00;
    end         
    
    endcase
end    
endmodule

